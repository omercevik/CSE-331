module muxLevel4(M, A, s4);
	input [31:0] A;
	input s4;
	output [31:0] M;
	
	mux2to1 m0(M[0], A[16], A[0], s4);
	mux2to1 m1(M[1], A[17], A[1], s4);
	mux2to1 m2(M[2], A[18], A[2], s4);
	mux2to1 m3(M[3], A[19], A[3], s4);
	mux2to1 m4(M[4], A[20], A[4], s4);
	mux2to1 m5(M[5], A[21], A[5], s4);
	mux2to1 m6(M[6], A[22], A[6], s4);
	mux2to1 m7(M[7], A[23], A[7], s4);
	mux2to1 m8(M[8], A[24], A[8], s4);
	mux2to1 m9(M[9], A[25], A[9], s4);
	mux2to1 m10(M[10], A[26], A[10], s4);
	mux2to1 m11(M[11], A[27], A[11], s4);
	mux2to1 m12(M[12], A[28], A[12], s4);
	mux2to1 m13(M[13], A[29], A[13], s4);
	mux2to1 m14(M[14], A[30], A[14], s4);
	mux2to1 m15(M[15], A[31], A[15], s4);
	mux2to1 m16(M[16], 1'b0, A[16], s4);
	mux2to1 m17(M[17], 1'b0, A[17], s4);
	mux2to1 m18(M[18], 1'b0, A[18], s4);
	mux2to1 m19(M[19], 1'b0, A[19], s4);
	mux2to1 m20(M[20], 1'b0, A[20], s4);
	mux2to1 m21(M[21], 1'b0, A[21], s4);
	mux2to1 m22(M[22], 1'b0, A[22], s4);
	mux2to1 m23(M[23], 1'b0, A[23], s4);
	mux2to1 m24(M[24], 1'b0, A[24], s4);
	mux2to1 m25(M[25], 1'b0, A[25], s4);
	mux2to1 m26(M[26], 1'b0, A[26], s4);
	mux2to1 m27(M[27], 1'b0, A[27], s4);
	mux2to1 m28(M[28], 1'b0, A[28], s4);
	mux2to1 m29(M[29], 1'b0, A[29], s4);
	mux2to1 m30(M[30], 1'b0, A[30], s4);
	mux2to1 m31(M[31], 1'b0, A[31], s4);
endmodule 