module orer(ored, a, b);
input [31:0]a, b;
output [31:0]ored;

or oring0(ored[0], a[0], b[0]);
or oring1(ored[1], a[1], b[1]);
or oring2(ored[2], a[2], b[2]);
or oring3(ored[3], a[3], b[3]);
or oring4(ored[4], a[4], b[4]);
or oring5(ored[5], a[5], b[5]);
or oring6(ored[6], a[6], b[6]);
or oring7(ored[7], a[7], b[7]);
or oring8(ored[8], a[8], b[8]);
or oring9(ored[9], a[9], b[9]);
or oring10(ored[10], a[10], b[10]);
or oring11(ored[11], a[11], b[11]);
or oring12(ored[12], a[12], b[12]);
or oring13(ored[13], a[13], b[13]);
or oring14(ored[14], a[14], b[14]);
or oring15(ored[15], a[15], b[15]);
or oring16(ored[16], a[16], b[16]);
or oring17(ored[17], a[17], b[17]);
or oring18(ored[18], a[18], b[18]);
or oring19(ored[19], a[19], b[19]);
or oring20(ored[20], a[20], b[20]);
or oring21(ored[21], a[21], b[21]);
or oring22(ored[22], a[22], b[22]);
or oring23(ored[23], a[23], b[23]);
or oring24(ored[24], a[24], b[24]);
or oring25(ored[25], a[25], b[25]);
or oring26(ored[26], a[26], b[26]);
or oring27(ored[27], a[27], b[27]);
or oring28(ored[28], a[28], b[28]);
or oring29(ored[29], a[29], b[29]);
or oring30(ored[30], a[30], b[30]);
or oring31(ored[31], a[31], b[31]);

endmodule 