module mips32_instruction_memory(read_address, instr);

	input [31:0] read_address;
	output [31:0] instr;
	
	
	initial
	begin
		
	end

	
	
endmodule 