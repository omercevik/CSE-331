module ander(anded, a, b);
input [31:0]a, b;
output [31:0]anded;

and anding0(anded[0], a[0], b[0]);
and anding1(anded[1], a[1], b[1]);
and anding2(anded[2], a[2], b[2]);
and anding3(anded[3], a[3], b[3]);
and anding4(anded[4], a[4], b[4]);
and anding5(anded[5], a[5], b[5]);
and anding6(anded[6], a[6], b[6]);
and anding7(anded[7], a[7], b[7]);
and anding8(anded[8], a[8], b[8]);
and anding9(anded[9], a[9], b[9]);
and anding10(anded[10], a[10], b[10]);
and anding11(anded[11], a[11], b[11]);
and anding12(anded[12], a[12], b[12]);
and anding13(anded[13], a[13], b[13]);
and anding14(anded[14], a[14], b[14]);
and anding15(anded[15], a[15], b[15]);
and anding16(anded[16], a[16], b[16]);
and anding17(anded[17], a[17], b[17]);
and anding18(anded[18], a[18], b[18]);
and anding19(anded[19], a[19], b[19]);
and anding20(anded[20], a[20], b[20]);
and anding21(anded[21], a[21], b[21]);
and anding22(anded[22], a[22], b[22]);
and anding23(anded[23], a[23], b[23]);
and anding24(anded[24], a[24], b[24]);
and anding25(anded[25], a[25], b[25]);
and anding26(anded[26], a[26], b[26]);
and anding27(anded[27], a[27], b[27]);
and anding28(anded[28], a[28], b[28]);
and anding29(anded[29], a[29], b[29]);
and anding30(anded[30], a[30], b[30]);
and anding31(anded[31], a[31], b[31]);

endmodule 