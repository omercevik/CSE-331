module norer(nored, a, b);
input [31:0]a, b;
output [31:0]nored;

nor noring0(nored[0], a[0], b[0]);
nor noring1(nored[1], a[1], b[1]);
nor noring2(nored[2], a[2], b[2]);
nor noring3(nored[3], a[3], b[3]);
nor noring4(nored[4], a[4], b[4]);
nor noring5(nored[5], a[5], b[5]);
nor noring6(nored[6], a[6], b[6]);
nor noring7(nored[7], a[7], b[7]);
nor noring8(nored[8], a[8], b[8]);
nor noring9(nored[9], a[9], b[9]);
nor noring10(nored[10], a[10], b[10]);
nor noring11(nored[11], a[11], b[11]);
nor noring12(nored[12], a[12], b[12]);
nor noring13(nored[13], a[13], b[13]);
nor noring14(nored[14], a[14], b[14]);
nor noring15(nored[15], a[15], b[15]);
nor noring16(nored[16], a[16], b[16]);
nor noring17(nored[17], a[17], b[17]);
nor noring18(nored[18], a[18], b[18]);
nor noring19(nored[19], a[19], b[19]);
nor noring20(nored[20], a[20], b[20]);
nor noring21(nored[21], a[21], b[21]);
nor noring22(nored[22], a[22], b[22]);
nor noring23(nored[23], a[23], b[23]);
nor noring24(nored[24], a[24], b[24]);
nor noring25(nored[25], a[25], b[25]);
nor noring26(nored[26], a[26], b[26]);
nor noring27(nored[27], a[27], b[27]);
nor noring28(nored[28], a[28], b[28]);
nor noring29(nored[29], a[29], b[29]);
nor noring30(nored[30], a[30], b[30]);
nor noring31(nored[31], a[31], b[31]);

endmodule 